/*   module top;

enum integer {a=0,b=5,c=7,d} var1;
initial
begin
$display(var1.first);
var1=b;
$display(var1.name);
var1=d;
$display(var1.prev);
$display(var1.num());
$display(var1.last); //8
end


endmodule       */



/* module top;

typedef enum time {a=1032,b=2003,c=2004,d=5000} t1;

t1 t2;
initial
begin
$display(t2.first);
t2=b;
$display(t2.name);
t2=d;
$display(t2.prev);
$display(t2.num());
$display(t2.last); 




end
endmodule */
